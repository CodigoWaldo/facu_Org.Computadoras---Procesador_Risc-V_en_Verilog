/*
Camino de datos: Conexiones que relacionan los distintos 
modulos para conformar el procesador.
*/


module datapath(
   
);


always @(*) 
    begin  
      
    end

endmodule